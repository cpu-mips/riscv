module asmtest(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h93031000;
30'h00000001: inst = 32'hb7000010;
30'h00000002: inst = 32'h93800002;
30'h00000003: inst = 32'h37b1ad1e;
30'h00000004: inst = 32'h1301f10e;
30'h00000005: inst = 32'h37050010;
30'h00000006: inst = 32'h23201500;
30'h00000007: inst = 32'h23222500;
30'h00000008: inst = 32'h83250500;
30'h00000009: inst = 32'h03264500;
30'h0000000a: inst = 32'h6394b014;
30'h0000000b: inst = 32'h93831300;
30'h0000000c: inst = 32'h6310c114;
30'h0000000d: inst = 32'h93831300;
30'h0000000e: inst = 32'h93831300;
30'h0000000f: inst = 32'h13048000;
30'h00000010: inst = 32'hb3047400;
30'h00000011: inst = 32'hb3a58400;
30'h00000012: inst = 32'h63940512;
30'h00000013: inst = 32'hb3259400;
30'h00000014: inst = 32'h63800512;
30'h00000015: inst = 32'h93a58400;
30'h00000016: inst = 32'h639c0510;
30'h00000017: inst = 32'h93831300;
30'h00000018: inst = 32'h13048000;
30'h00000019: inst = 32'h93543400;
30'h0000001a: inst = 32'h93051000;
30'h0000001b: inst = 32'h6392b410;
30'h0000001c: inst = 32'hb394b400;
30'h0000001d: inst = 32'h13062000;
30'h0000001e: inst = 32'h631c960e;
30'h0000001f: inst = 32'h93831300;
30'h00000020: inst = 32'h9304f000;
30'h00000021: inst = 32'hb3e50400;
30'h00000022: inst = 32'h6394b40e;
30'h00000023: inst = 32'hb3c50400;
30'h00000024: inst = 32'h6390950e;
30'h00000025: inst = 32'hb3f50400;
30'h00000026: inst = 32'h639c050c;
30'h00000027: inst = 32'h93831300;
30'h00000028: inst = 32'h83250500;
30'h00000029: inst = 32'hb384a500;
30'h0000002a: inst = 32'h93858500;
30'h0000002b: inst = 32'h23a09500;
30'h0000002c: inst = 32'h03a60500;
30'h0000002d: inst = 32'h639ec40a;
30'h0000002e: inst = 32'h13000000;
30'h0000002f: inst = 32'h93831300;
30'h00000030: inst = 32'h93040000;
30'h00000031: inst = 32'h6f004000;
30'h00000032: inst = 32'h13040000;
30'h00000033: inst = 32'h6312940a;
30'h00000034: inst = 32'h33808300;
30'h00000035: inst = 32'h631e8008;
30'h00000036: inst = 32'h93850300;
30'h00000037: inst = 32'h93831300;
30'h00000038: inst = 32'h63887508;
30'h00000039: inst = 32'h63c6b308;
30'h0000003a: inst = 32'h63c47308;
30'h0000003b: inst = 32'h63d27508;
30'h0000003c: inst = 32'h63907308;
30'h0000003d: inst = 32'h37f4ffff;
30'h0000003e: inst = 32'h13041400;
30'h0000003f: inst = 32'h37010000;
30'h00000040: inst = 32'h13011100;
30'h00000041: inst = 32'h63662406;
30'h00000042: inst = 32'h63648406;
30'h00000043: inst = 32'h63728106;
30'h00000044: inst = 32'h93831300;
30'h00000045: inst = 32'h37b4adde;
30'h00000046: inst = 32'h1304f40e;
30'h00000047: inst = 32'h9300f00e;
30'h00000048: inst = 32'h37b10000;
30'h00000049: inst = 32'h1301f10e;
30'h0000004a: inst = 32'hb7f1ffff;
30'h0000004b: inst = 32'h9302f000;
30'h0000004c: inst = 32'h93928200;
30'h0000004d: inst = 32'hb3813200;
30'h0000004e: inst = 32'h9381f10e;
30'h0000004f: inst = 32'h37b2ffff;
30'h00000050: inst = 32'h1302f20e;
30'h00000051: inst = 32'h23008502;
30'h00000052: inst = 32'h23108504;
30'h00000053: inst = 32'h83440502;
30'h00000054: inst = 32'h83550504;
30'h00000055: inst = 32'h83020502;
30'h00000056: inst = 32'h03130504;
30'h00000057: inst = 32'h639a1400;
30'h00000058: inst = 32'h63982500;
30'h00000059: inst = 32'h63963200;
30'h0000005a: inst = 32'h63144300;
30'h0000005b: inst = 32'h6f008004;
30'h0000005c: inst = 32'h13026004;
30'h0000005d: inst = 32'hef000007;
30'h0000005e: inst = 32'h13021006;
30'h0000005f: inst = 32'hef008006;
30'h00000060: inst = 32'h13029006;
30'h00000061: inst = 32'hef000006;
30'h00000062: inst = 32'h1302c006;
30'h00000063: inst = 32'hef008005;
30'h00000064: inst = 32'h1302a003;
30'h00000065: inst = 32'hef000005;
30'h00000066: inst = 32'h13020002;
30'h00000067: inst = 32'hef008004;
30'h00000068: inst = 32'h13820303;
30'h00000069: inst = 32'hef000004;
30'h0000006a: inst = 32'h1302a000;
30'h0000006b: inst = 32'hef008003;
30'h0000006c: inst = 32'h6f000003;
30'h0000006d: inst = 32'h13020005;
30'h0000006e: inst = 32'hef00c002;
30'h0000006f: inst = 32'h13021006;
30'h00000070: inst = 32'hef004002;
30'h00000071: inst = 32'h13023007;
30'h00000072: inst = 32'hef00c001;
30'h00000073: inst = 32'h13023007;
30'h00000074: inst = 32'hef004001;
30'h00000075: inst = 32'h1302a000;
30'h00000076: inst = 32'hef00c000;
30'h00000077: inst = 32'h6f004000;
30'h00000078: inst = 32'h6f000000;
30'h00000079: inst = 32'h37010080;
30'h0000007a: inst = 32'h83210100;
30'h0000007b: inst = 32'h93f11100;
30'h0000007c: inst = 32'he38a01fe;
30'h0000007d: inst = 32'h23244100;
30'h0000007e: inst = 32'h67800000;
default:      inst = 32'h00000000;
endcase
end
endmodule
