module example(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h37070010;
30'h00000001: inst = 32'h13070760;
30'h00000002: inst = 32'hef004000;
30'h00000003: inst = 32'h130707fd;
30'h00000004: inst = 32'h23262702;
30'h00000005: inst = 32'h13010703;
30'h00000006: inst = 32'h13084006;
30'h00000007: inst = 32'h232601ff;
30'h00000008: inst = 32'h0328c1fe;
30'h00000009: inst = 32'h1308481f;
30'h0000000a: inst = 32'h232401ff;
30'h0000000b: inst = 32'h1308803e;
30'h0000000c: inst = 32'h232201ff;
30'h0000000d: inst = 32'h032841fe;
30'h0000000e: inst = 32'h1348f8ff;
30'h0000000f: inst = 32'h232001ff;
30'h00000010: inst = 32'h37080010;
30'h00000011: inst = 32'h1308880f;
30'h00000012: inst = 32'h03483800;
30'h00000013: inst = 32'ha30f01fd;
30'h00000014: inst = 32'h37080010;
30'h00000015: inst = 32'h1308880f;
30'h00000016: inst = 32'h93082004;
30'h00000017: inst = 32'h23021801;
30'h00000018: inst = 32'h37080010;
30'h00000019: inst = 32'h1308880f;
30'h0000001a: inst = 32'h93083004;
30'h0000001b: inst = 32'ha3021801;
30'h0000001c: inst = 32'h37080010;
30'h0000001d: inst = 32'h1308880f;
30'h0000001e: inst = 32'h93084004;
30'h0000001f: inst = 32'h23031801;
30'h00000020: inst = 32'h37080010;
30'h00000021: inst = 32'h1308880f;
30'h00000022: inst = 32'h93085004;
30'h00000023: inst = 32'ha3031801;
30'h00000024: inst = 32'h37080010;
30'h00000025: inst = 32'h1308880f;
30'h00000026: inst = 32'h03484800;
30'h00000027: inst = 32'h230f01fd;
30'h00000028: inst = 32'h37080010;
30'h00000029: inst = 32'h1308880f;
30'h0000002a: inst = 32'h03485800;
30'h0000002b: inst = 32'ha30e01fd;
30'h0000002c: inst = 32'h37080010;
30'h0000002d: inst = 32'h1308880f;
30'h0000002e: inst = 32'h03486800;
30'h0000002f: inst = 32'h230e01fd;
30'h00000030: inst = 32'h37080010;
30'h00000031: inst = 32'h1308880f;
30'h00000032: inst = 32'h03487800;
30'h00000033: inst = 32'ha30d01fd;
30'h00000034: inst = 32'h032881fe;
30'h00000035: inst = 32'h0321c702;
30'h00000036: inst = 32'h13070703;
30'h00000037: inst = 32'h67800000;
30'h00000038: inst = 32'h03000000;
30'h00000039: inst = 32'h02000000;
30'h0000003a: inst = 32'h04000000;
30'h0000003b: inst = 32'h17000000;
30'h0000003c: inst = 32'h20000000;
30'h0000003d: inst = 32'h01000000;
30'h0000003e: inst = 32'h48454c4c;
30'h0000003f: inst = 32'h4f20574f;
30'h00000040: inst = 32'h524c4421;
30'h00000041: inst = 32'h21000000;
default:      inst = 32'h00000000;
endcase
end
endmodule
